module core();
endmodule